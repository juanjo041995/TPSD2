----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:34:28 10/16/2020 
-- Design Name: 
-- Module Name:    PruebaDualRam - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity PruebaDualRam is
	PORT (
				clk : in STD_LOGIC;
				reset: in STD_LOGIC;
				HSync: out STD_LOGIC;
				
	);
end PruebaDualRam;

architecture Behavioral of PruebaDualRam is

begin


end Behavioral;

