----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:55:34 10/20/2020 
-- Design Name: 
-- Module Name:    pauseIn - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity pauseIn is
	PORT (
				SW3,SW4 : in STD_LOGIC;
				clk	  : in STD_LOGIC;
				pause	  : out STD_LOGIC :='0'
	);
end pauseIn;

architecture Behavioral of pauseIn is

begin
		process (clk)
		begin
			if (clk'event and clk='1') then
				if SW4 = '0' then
					pause <= '1';
				elsif SW3 = '0' then
					pause <= '0';
				end if;
			end if;
		end process;

end Behavioral;

